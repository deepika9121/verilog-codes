`timescale 1ns / 1ps
// Engineer: B DEEPIKA
// Design Name: fulladder using demux1x8
// Module Name: fulladder_using_demux1x8
/////////////////////////////////////////


module fulladder_using_demux1x8();

endmodule
